module rw_control_logic(dataBuffer,groupControl,portControl,RD_bar,WR_bar,
A0,A1,CS_bar,RESET);

output dataBuffer, groupControl, portControl;
//dataBuffer => output from control logic to data buffer 
//groupControl => output from control logic to group A&B control 
//portControl => output from control logic to port A,B&C 

input RD_bar, WR_bar, A0, A1, CS_bar, RESET;
//RD_bar => read data from ports to CPU
//WR_bar => write data from CPU to Ports
//A0 & A1 => Port selection
//CS_bar => enable of chip
//RESET => reset signal











endmodule

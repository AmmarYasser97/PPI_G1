module INOUT_mode(DATA, A0, A1);
input [7:0]Control;



endmodule
